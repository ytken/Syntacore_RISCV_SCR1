// de10lite_sopc.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module de10lite_sopc (
		output wire        avl_dmem_waitrequest,   //        avl_dmem.waitrequest
		output wire [31:0] avl_dmem_readdata,      //                .readdata
		output wire        avl_dmem_readdatavalid, //                .readdatavalid
		output wire [1:0]  avl_dmem_response,      //                .response
		input  wire [0:0]  avl_dmem_burstcount,    //                .burstcount
		input  wire [31:0] avl_dmem_writedata,     //                .writedata
		input  wire [31:0] avl_dmem_address,       //                .address
		input  wire        avl_dmem_write,         //                .write
		input  wire        avl_dmem_read,          //                .read
		input  wire [3:0]  avl_dmem_byteenable,    //                .byteenable
		input  wire        avl_dmem_debugaccess,   //                .debugaccess
		output wire        avl_imem_waitrequest,   //        avl_imem.waitrequest
		output wire [31:0] avl_imem_readdata,      //                .readdata
		output wire        avl_imem_readdatavalid, //                .readdatavalid
		output wire [1:0]  avl_imem_response,      //                .response
		input  wire [0:0]  avl_imem_burstcount,    //                .burstcount
		input  wire [31:0] avl_imem_writedata,     //                .writedata
		input  wire [31:0] avl_imem_address,       //                .address
		input  wire        avl_imem_write,         //                .write
		input  wire        avl_imem_read,          //                .read
		input  wire [3:0]  avl_imem_byteenable,    //                .byteenable
		input  wire        avl_imem_debugaccess,   //                .debugaccess
		input  wire [31:0] bld_id_export,          //          bld_id.export
		input  wire [31:0] core_clk_freq_export,   //   core_clk_freq.export
		output wire        cpu_clk_out_clk,        //     cpu_clk_out.clk
		output wire        cpu_rst_out_reset_n,    //     cpu_rst_out.reset_n
		input  wire        osc_50_clk,             //          osc_50.clk
		output wire [18:0] pio_led_export,         //         pio_led.export
		input  wire [18:0] pio_sw_export,          //          pio_sw.export
		input  wire        pll_reset,              //             pll.reset
		output wire        pwrup_rst_n_out_export, // pwrup_rst_n_out.export
		output wire [12:0] sdram_addr,             //           sdram.addr
		output wire [1:0]  sdram_ba,               //                .ba
		output wire        sdram_cas_n,            //                .cas_n
		output wire        sdram_cke,              //                .cke
		output wire        sdram_cs_n,             //                .cs_n
		inout  wire [15:0] sdram_dq,               //                .dq
		output wire [1:0]  sdram_dqm,              //                .dqm
		output wire        sdram_ras_n,            //                .ras_n
		output wire        sdram_we_n,             //                .we_n
		output wire        sdram_clk_out_clk,      //   sdram_clk_out.clk
		input  wire        soc_reset_n,            //             soc.reset_n
		input  wire [31:0] soc_id_export,          //          soc_id.export
		input  wire        uart_waitrequest,       //            uart.waitrequest
		input  wire [31:0] uart_readdata,          //                .readdata
		input  wire        uart_readdatavalid,     //                .readdatavalid
		output wire [0:0]  uart_burstcount,        //                .burstcount
		output wire [31:0] uart_writedata,         //                .writedata
		output wire [4:0]  uart_address,           //                .address
		output wire        uart_write,             //                .write
		output wire        uart_read,              //                .read
		output wire [3:0]  uart_byteenable,        //                .byteenable
		output wire        uart_debugaccess        //                .debugaccess
	);

	wire         pll_0_outclk1_clk;                                    // pll_0:outclk_1 -> [mm_interconnect_0:pll_0_outclk1_clk, rst_controller_002:clk, sdram:clk]
	wire         avl_imem_m0_waitrequest;                              // mm_interconnect_0:avl_imem_m0_waitrequest -> avl_imem:m0_waitrequest
	wire  [31:0] avl_imem_m0_readdata;                                 // mm_interconnect_0:avl_imem_m0_readdata -> avl_imem:m0_readdata
	wire         avl_imem_m0_debugaccess;                              // avl_imem:m0_debugaccess -> mm_interconnect_0:avl_imem_m0_debugaccess
	wire  [31:0] avl_imem_m0_address;                                  // avl_imem:m0_address -> mm_interconnect_0:avl_imem_m0_address
	wire         avl_imem_m0_read;                                     // avl_imem:m0_read -> mm_interconnect_0:avl_imem_m0_read
	wire   [3:0] avl_imem_m0_byteenable;                               // avl_imem:m0_byteenable -> mm_interconnect_0:avl_imem_m0_byteenable
	wire         avl_imem_m0_readdatavalid;                            // mm_interconnect_0:avl_imem_m0_readdatavalid -> avl_imem:m0_readdatavalid
	wire   [1:0] avl_imem_m0_response;                                 // mm_interconnect_0:avl_imem_m0_response -> avl_imem:m0_response
	wire  [31:0] avl_imem_m0_writedata;                                // avl_imem:m0_writedata -> mm_interconnect_0:avl_imem_m0_writedata
	wire         avl_imem_m0_write;                                    // avl_imem:m0_write -> mm_interconnect_0:avl_imem_m0_write
	wire   [0:0] avl_imem_m0_burstcount;                               // avl_imem:m0_burstcount -> mm_interconnect_0:avl_imem_m0_burstcount
	wire         avl_dmem_m0_waitrequest;                              // mm_interconnect_0:avl_dmem_m0_waitrequest -> avl_dmem:m0_waitrequest
	wire  [31:0] avl_dmem_m0_readdata;                                 // mm_interconnect_0:avl_dmem_m0_readdata -> avl_dmem:m0_readdata
	wire         avl_dmem_m0_debugaccess;                              // avl_dmem:m0_debugaccess -> mm_interconnect_0:avl_dmem_m0_debugaccess
	wire  [31:0] avl_dmem_m0_address;                                  // avl_dmem:m0_address -> mm_interconnect_0:avl_dmem_m0_address
	wire         avl_dmem_m0_read;                                     // avl_dmem:m0_read -> mm_interconnect_0:avl_dmem_m0_read
	wire   [3:0] avl_dmem_m0_byteenable;                               // avl_dmem:m0_byteenable -> mm_interconnect_0:avl_dmem_m0_byteenable
	wire         avl_dmem_m0_readdatavalid;                            // mm_interconnect_0:avl_dmem_m0_readdatavalid -> avl_dmem:m0_readdatavalid
	wire   [1:0] avl_dmem_m0_response;                                 // mm_interconnect_0:avl_dmem_m0_response -> avl_dmem:m0_response
	wire  [31:0] avl_dmem_m0_writedata;                                // avl_dmem:m0_writedata -> mm_interconnect_0:avl_dmem_m0_writedata
	wire         avl_dmem_m0_write;                                    // avl_dmem:m0_write -> mm_interconnect_0:avl_dmem_m0_write
	wire   [0:0] avl_dmem_m0_burstcount;                               // avl_dmem:m0_burstcount -> mm_interconnect_0:avl_dmem_m0_burstcount
	wire   [1:0] mm_interconnect_0_default_slave_axi_error_if_awburst; // mm_interconnect_0:default_slave_axi_error_if_awburst -> default_slave:awburst
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_arlen;   // mm_interconnect_0:default_slave_axi_error_if_arlen -> default_slave:arlen
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_wstrb;   // mm_interconnect_0:default_slave_axi_error_if_wstrb -> default_slave:wstrb
	wire         mm_interconnect_0_default_slave_axi_error_if_wready;  // default_slave:wready -> mm_interconnect_0:default_slave_axi_error_if_wready
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_rid;     // default_slave:rid -> mm_interconnect_0:default_slave_axi_error_if_rid
	wire         mm_interconnect_0_default_slave_axi_error_if_rready;  // mm_interconnect_0:default_slave_axi_error_if_rready -> default_slave:rready
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_awlen;   // mm_interconnect_0:default_slave_axi_error_if_awlen -> default_slave:awlen
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_wid;     // mm_interconnect_0:default_slave_axi_error_if_wid -> default_slave:wid
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_arcache; // mm_interconnect_0:default_slave_axi_error_if_arcache -> default_slave:arcache
	wire         mm_interconnect_0_default_slave_axi_error_if_wvalid;  // mm_interconnect_0:default_slave_axi_error_if_wvalid -> default_slave:wvalid
	wire  [31:0] mm_interconnect_0_default_slave_axi_error_if_araddr;  // mm_interconnect_0:default_slave_axi_error_if_araddr -> default_slave:araddr
	wire   [2:0] mm_interconnect_0_default_slave_axi_error_if_arprot;  // mm_interconnect_0:default_slave_axi_error_if_arprot -> default_slave:arprot
	wire   [2:0] mm_interconnect_0_default_slave_axi_error_if_awprot;  // mm_interconnect_0:default_slave_axi_error_if_awprot -> default_slave:awprot
	wire  [31:0] mm_interconnect_0_default_slave_axi_error_if_wdata;   // mm_interconnect_0:default_slave_axi_error_if_wdata -> default_slave:wdata
	wire         mm_interconnect_0_default_slave_axi_error_if_arvalid; // mm_interconnect_0:default_slave_axi_error_if_arvalid -> default_slave:arvalid
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_awcache; // mm_interconnect_0:default_slave_axi_error_if_awcache -> default_slave:awcache
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_arid;    // mm_interconnect_0:default_slave_axi_error_if_arid -> default_slave:arid
	wire   [1:0] mm_interconnect_0_default_slave_axi_error_if_arlock;  // mm_interconnect_0:default_slave_axi_error_if_arlock -> default_slave:arlock
	wire   [1:0] mm_interconnect_0_default_slave_axi_error_if_awlock;  // mm_interconnect_0:default_slave_axi_error_if_awlock -> default_slave:awlock
	wire  [31:0] mm_interconnect_0_default_slave_axi_error_if_awaddr;  // mm_interconnect_0:default_slave_axi_error_if_awaddr -> default_slave:awaddr
	wire   [1:0] mm_interconnect_0_default_slave_axi_error_if_bresp;   // default_slave:bresp -> mm_interconnect_0:default_slave_axi_error_if_bresp
	wire         mm_interconnect_0_default_slave_axi_error_if_arready; // default_slave:arready -> mm_interconnect_0:default_slave_axi_error_if_arready
	wire  [31:0] mm_interconnect_0_default_slave_axi_error_if_rdata;   // default_slave:rdata -> mm_interconnect_0:default_slave_axi_error_if_rdata
	wire         mm_interconnect_0_default_slave_axi_error_if_awready; // default_slave:awready -> mm_interconnect_0:default_slave_axi_error_if_awready
	wire   [1:0] mm_interconnect_0_default_slave_axi_error_if_arburst; // mm_interconnect_0:default_slave_axi_error_if_arburst -> default_slave:arburst
	wire   [2:0] mm_interconnect_0_default_slave_axi_error_if_arsize;  // mm_interconnect_0:default_slave_axi_error_if_arsize -> default_slave:arsize
	wire         mm_interconnect_0_default_slave_axi_error_if_bready;  // mm_interconnect_0:default_slave_axi_error_if_bready -> default_slave:bready
	wire         mm_interconnect_0_default_slave_axi_error_if_rlast;   // default_slave:rlast -> mm_interconnect_0:default_slave_axi_error_if_rlast
	wire         mm_interconnect_0_default_slave_axi_error_if_wlast;   // mm_interconnect_0:default_slave_axi_error_if_wlast -> default_slave:wlast
	wire   [1:0] mm_interconnect_0_default_slave_axi_error_if_rresp;   // default_slave:rresp -> mm_interconnect_0:default_slave_axi_error_if_rresp
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_awid;    // mm_interconnect_0:default_slave_axi_error_if_awid -> default_slave:awid
	wire   [3:0] mm_interconnect_0_default_slave_axi_error_if_bid;     // default_slave:bid -> mm_interconnect_0:default_slave_axi_error_if_bid
	wire         mm_interconnect_0_default_slave_axi_error_if_bvalid;  // default_slave:bvalid -> mm_interconnect_0:default_slave_axi_error_if_bvalid
	wire   [2:0] mm_interconnect_0_default_slave_axi_error_if_awsize;  // mm_interconnect_0:default_slave_axi_error_if_awsize -> default_slave:awsize
	wire         mm_interconnect_0_default_slave_axi_error_if_awvalid; // mm_interconnect_0:default_slave_axi_error_if_awvalid -> default_slave:awvalid
	wire         mm_interconnect_0_default_slave_axi_error_if_rvalid;  // default_slave:rvalid -> mm_interconnect_0:default_slave_axi_error_if_rvalid
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;           // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [63:0] mm_interconnect_0_onchip_ram_s1_readdata;             // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_ram_s1_address;              // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [7:0] mm_interconnect_0_onchip_ram_s1_byteenable;           // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [63:0] mm_interconnect_0_onchip_ram_s1_writedata;            // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                  // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;               // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                   // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                      // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;             // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                     // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                 // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_avl_uart_s0_readdata;               // avl_uart:s0_readdata -> mm_interconnect_0:avl_uart_s0_readdata
	wire         mm_interconnect_0_avl_uart_s0_waitrequest;            // avl_uart:s0_waitrequest -> mm_interconnect_0:avl_uart_s0_waitrequest
	wire         mm_interconnect_0_avl_uart_s0_debugaccess;            // mm_interconnect_0:avl_uart_s0_debugaccess -> avl_uart:s0_debugaccess
	wire   [4:0] mm_interconnect_0_avl_uart_s0_address;                // mm_interconnect_0:avl_uart_s0_address -> avl_uart:s0_address
	wire         mm_interconnect_0_avl_uart_s0_read;                   // mm_interconnect_0:avl_uart_s0_read -> avl_uart:s0_read
	wire   [3:0] mm_interconnect_0_avl_uart_s0_byteenable;             // mm_interconnect_0:avl_uart_s0_byteenable -> avl_uart:s0_byteenable
	wire         mm_interconnect_0_avl_uart_s0_readdatavalid;          // avl_uart:s0_readdatavalid -> mm_interconnect_0:avl_uart_s0_readdatavalid
	wire         mm_interconnect_0_avl_uart_s0_write;                  // mm_interconnect_0:avl_uart_s0_write -> avl_uart:s0_write
	wire  [31:0] mm_interconnect_0_avl_uart_s0_writedata;              // mm_interconnect_0:avl_uart_s0_writedata -> avl_uart:s0_writedata
	wire   [0:0] mm_interconnect_0_avl_uart_s0_burstcount;             // mm_interconnect_0:avl_uart_s0_burstcount -> avl_uart:s0_burstcount
	wire         mm_interconnect_0_pio_led_s1_chipselect;              // mm_interconnect_0:pio_led_s1_chipselect -> pio_led:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_s1_readdata;                // pio_led:readdata -> mm_interconnect_0:pio_led_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_led_s1_address;                 // mm_interconnect_0:pio_led_s1_address -> pio_led:address
	wire         mm_interconnect_0_pio_led_s1_write;                   // mm_interconnect_0:pio_led_s1_write -> pio_led:write_n
	wire  [31:0] mm_interconnect_0_pio_led_s1_writedata;               // mm_interconnect_0:pio_led_s1_writedata -> pio_led:writedata
	wire  [31:0] mm_interconnect_0_pio_sw_s1_readdata;                 // pio_sw:readdata -> mm_interconnect_0:pio_sw_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_sw_s1_address;                  // mm_interconnect_0:pio_sw_s1_address -> pio_sw:address
	wire  [31:0] mm_interconnect_0_bld_id_s1_readdata;                 // bld_id:readdata -> mm_interconnect_0:bld_id_s1_readdata
	wire   [1:0] mm_interconnect_0_bld_id_s1_address;                  // mm_interconnect_0:bld_id_s1_address -> bld_id:address
	wire  [31:0] mm_interconnect_0_soc_id_s1_readdata;                 // soc_id:readdata -> mm_interconnect_0:soc_id_s1_readdata
	wire   [1:0] mm_interconnect_0_soc_id_s1_address;                  // mm_interconnect_0:soc_id_s1_address -> soc_id:address
	wire  [31:0] mm_interconnect_0_core_clk_freq_s1_readdata;          // core_clk_freq:readdata -> mm_interconnect_0:core_clk_freq_s1_readdata
	wire   [1:0] mm_interconnect_0_core_clk_freq_s1_address;           // mm_interconnect_0:core_clk_freq_s1_address -> core_clk_freq:address
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [avl_dmem:reset, avl_imem:reset, avl_uart:reset, bld_id:reset_n, core_clk_freq:reset_n, default_slave:aresetn, mm_interconnect_0:avl_imem_reset_reset_bridge_in_reset_reset, onchip_ram:reset, pio_led:reset_n, pio_sw:reset_n, soc_id:reset_n]
	wire         reset_sequencer_0_reset_out0_reset;                   // reset_sequencer_0:reset_out0 -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	wire         rst_controller_001_reset_out_reset;                   // rst_controller_001:reset_out -> rst_controller_001_reset_out_reset:in
	wire         reset_sequencer_0_reset_out1_reset;                   // reset_sequencer_0:reset_out1 -> rst_controller_001:reset_in0
	wire         rst_controller_002_reset_out_reset;                   // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, sdram:reset_n]

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) avl_dmem (
		.clk              (cpu_clk_out_clk),                //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (avl_dmem_waitrequest),           //    s0.waitrequest
		.s0_readdata      (avl_dmem_readdata),              //      .readdata
		.s0_readdatavalid (avl_dmem_readdatavalid),         //      .readdatavalid
		.s0_response      (avl_dmem_response),              //      .response
		.s0_burstcount    (avl_dmem_burstcount),            //      .burstcount
		.s0_writedata     (avl_dmem_writedata),             //      .writedata
		.s0_address       (avl_dmem_address),               //      .address
		.s0_write         (avl_dmem_write),                 //      .write
		.s0_read          (avl_dmem_read),                  //      .read
		.s0_byteenable    (avl_dmem_byteenable),            //      .byteenable
		.s0_debugaccess   (avl_dmem_debugaccess),           //      .debugaccess
		.m0_waitrequest   (avl_dmem_m0_waitrequest),        //    m0.waitrequest
		.m0_readdata      (avl_dmem_m0_readdata),           //      .readdata
		.m0_readdatavalid (avl_dmem_m0_readdatavalid),      //      .readdatavalid
		.m0_response      (avl_dmem_m0_response),           //      .response
		.m0_burstcount    (avl_dmem_m0_burstcount),         //      .burstcount
		.m0_writedata     (avl_dmem_m0_writedata),          //      .writedata
		.m0_address       (avl_dmem_m0_address),            //      .address
		.m0_write         (avl_dmem_m0_write),              //      .write
		.m0_read          (avl_dmem_m0_read),               //      .read
		.m0_byteenable    (avl_dmem_m0_byteenable),         //      .byteenable
		.m0_debugaccess   (avl_dmem_m0_debugaccess)         //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) avl_imem (
		.clk              (cpu_clk_out_clk),                //   clk.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.s0_waitrequest   (avl_imem_waitrequest),           //    s0.waitrequest
		.s0_readdata      (avl_imem_readdata),              //      .readdata
		.s0_readdatavalid (avl_imem_readdatavalid),         //      .readdatavalid
		.s0_response      (avl_imem_response),              //      .response
		.s0_burstcount    (avl_imem_burstcount),            //      .burstcount
		.s0_writedata     (avl_imem_writedata),             //      .writedata
		.s0_address       (avl_imem_address),               //      .address
		.s0_write         (avl_imem_write),                 //      .write
		.s0_read          (avl_imem_read),                  //      .read
		.s0_byteenable    (avl_imem_byteenable),            //      .byteenable
		.s0_debugaccess   (avl_imem_debugaccess),           //      .debugaccess
		.m0_waitrequest   (avl_imem_m0_waitrequest),        //    m0.waitrequest
		.m0_readdata      (avl_imem_m0_readdata),           //      .readdata
		.m0_readdatavalid (avl_imem_m0_readdatavalid),      //      .readdatavalid
		.m0_response      (avl_imem_m0_response),           //      .response
		.m0_burstcount    (avl_imem_m0_burstcount),         //      .burstcount
		.m0_writedata     (avl_imem_m0_writedata),          //      .writedata
		.m0_address       (avl_imem_m0_address),            //      .address
		.m0_write         (avl_imem_m0_write),              //      .write
		.m0_read          (avl_imem_m0_read),               //      .read
		.m0_byteenable    (avl_imem_m0_byteenable),         //      .byteenable
		.m0_debugaccess   (avl_imem_m0_debugaccess)         //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (5),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) avl_uart (
		.clk              (cpu_clk_out_clk),                             //   clk.clk
		.reset            (rst_controller_reset_out_reset),              // reset.reset
		.s0_waitrequest   (mm_interconnect_0_avl_uart_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_avl_uart_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_avl_uart_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_avl_uart_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_avl_uart_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_avl_uart_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_avl_uart_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_avl_uart_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_avl_uart_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_avl_uart_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (uart_waitrequest),                            //    m0.waitrequest
		.m0_readdata      (uart_readdata),                               //      .readdata
		.m0_readdatavalid (uart_readdatavalid),                          //      .readdatavalid
		.m0_burstcount    (uart_burstcount),                             //      .burstcount
		.m0_writedata     (uart_writedata),                              //      .writedata
		.m0_address       (uart_address),                                //      .address
		.m0_write         (uart_write),                                  //      .write
		.m0_read          (uart_read),                                   //      .read
		.m0_byteenable    (uart_byteenable),                             //      .byteenable
		.m0_debugaccess   (uart_debugaccess),                            //      .debugaccess
		.s0_response      (),                                            // (terminated)
		.m0_response      (2'b00)                                        // (terminated)
	);

	de10lite_sopc_bld_id bld_id (
		.clk      (cpu_clk_out_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_bld_id_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_bld_id_s1_readdata), //                    .readdata
		.in_port  (bld_id_export)                         // external_connection.export
	);

	de10lite_sopc_core_clk_freq core_clk_freq (
		.clk      (cpu_clk_out_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_core_clk_freq_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_core_clk_freq_s1_readdata), //                    .readdata
		.in_port  (core_clk_freq_export)                         // external_connection.export
	);

	altera_error_response_slave #(
		.AXI_ID_W           (4),
		.AXI_ADDR_W         (32),
		.AXI_DATA_W         (32),
		.SUPPORT_CSR        (0),
		.LOG_CSR_DEPTH      (1),
		.REGISTER_AV_INPUTS (0)
	) default_slave (
		.aclk    (cpu_clk_out_clk),                                      //          clk.clk
		.aresetn (~rst_controller_reset_out_reset),                      //    clk_reset.reset_n
		.awid    (mm_interconnect_0_default_slave_axi_error_if_awid),    // axi_error_if.awid
		.awaddr  (mm_interconnect_0_default_slave_axi_error_if_awaddr),  //             .awaddr
		.awlen   (mm_interconnect_0_default_slave_axi_error_if_awlen),   //             .awlen
		.awsize  (mm_interconnect_0_default_slave_axi_error_if_awsize),  //             .awsize
		.awburst (mm_interconnect_0_default_slave_axi_error_if_awburst), //             .awburst
		.awlock  (mm_interconnect_0_default_slave_axi_error_if_awlock),  //             .awlock
		.awcache (mm_interconnect_0_default_slave_axi_error_if_awcache), //             .awcache
		.awprot  (mm_interconnect_0_default_slave_axi_error_if_awprot),  //             .awprot
		.awvalid (mm_interconnect_0_default_slave_axi_error_if_awvalid), //             .awvalid
		.awready (mm_interconnect_0_default_slave_axi_error_if_awready), //             .awready
		.wid     (mm_interconnect_0_default_slave_axi_error_if_wid),     //             .wid
		.wdata   (mm_interconnect_0_default_slave_axi_error_if_wdata),   //             .wdata
		.wstrb   (mm_interconnect_0_default_slave_axi_error_if_wstrb),   //             .wstrb
		.wlast   (mm_interconnect_0_default_slave_axi_error_if_wlast),   //             .wlast
		.wvalid  (mm_interconnect_0_default_slave_axi_error_if_wvalid),  //             .wvalid
		.wready  (mm_interconnect_0_default_slave_axi_error_if_wready),  //             .wready
		.bid     (mm_interconnect_0_default_slave_axi_error_if_bid),     //             .bid
		.bresp   (mm_interconnect_0_default_slave_axi_error_if_bresp),   //             .bresp
		.bvalid  (mm_interconnect_0_default_slave_axi_error_if_bvalid),  //             .bvalid
		.bready  (mm_interconnect_0_default_slave_axi_error_if_bready),  //             .bready
		.arid    (mm_interconnect_0_default_slave_axi_error_if_arid),    //             .arid
		.araddr  (mm_interconnect_0_default_slave_axi_error_if_araddr),  //             .araddr
		.arlen   (mm_interconnect_0_default_slave_axi_error_if_arlen),   //             .arlen
		.arsize  (mm_interconnect_0_default_slave_axi_error_if_arsize),  //             .arsize
		.arburst (mm_interconnect_0_default_slave_axi_error_if_arburst), //             .arburst
		.arlock  (mm_interconnect_0_default_slave_axi_error_if_arlock),  //             .arlock
		.arcache (mm_interconnect_0_default_slave_axi_error_if_arcache), //             .arcache
		.arprot  (mm_interconnect_0_default_slave_axi_error_if_arprot),  //             .arprot
		.arvalid (mm_interconnect_0_default_slave_axi_error_if_arvalid), //             .arvalid
		.arready (mm_interconnect_0_default_slave_axi_error_if_arready), //             .arready
		.rid     (mm_interconnect_0_default_slave_axi_error_if_rid),     //             .rid
		.rdata   (mm_interconnect_0_default_slave_axi_error_if_rdata),   //             .rdata
		.rresp   (mm_interconnect_0_default_slave_axi_error_if_rresp),   //             .rresp
		.rlast   (mm_interconnect_0_default_slave_axi_error_if_rlast),   //             .rlast
		.rvalid  (mm_interconnect_0_default_slave_axi_error_if_rvalid),  //             .rvalid
		.rready  (mm_interconnect_0_default_slave_axi_error_if_rready)   //             .rready
	);

	de10lite_sopc_onchip_ram onchip_ram (
		.clk        (cpu_clk_out_clk),                            //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (1'b0),                                       // (terminated)
		.freeze     (1'b0)                                        // (terminated)
	);

	de10lite_sopc_pio_led pio_led (
		.clk        (cpu_clk_out_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_export)                           // external_connection.export
	);

	de10lite_sopc_pio_sw pio_sw (
		.clk      (cpu_clk_out_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_pio_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_sw_s1_readdata), //                    .readdata
		.in_port  (pio_sw_export)                         // external_connection.export
	);

	de10lite_sopc_pll_0 pll_0 (
		.refclk   (osc_50_clk),             //  refclk.clk
		.rst      (pll_reset),              //   reset.reset
		.outclk_0 (cpu_clk_out_clk),        // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk),      // outclk1.clk
		.outclk_2 (sdram_clk_out_clk),      // outclk2.clk
		.locked   (pwrup_rst_n_out_export)  //  locked.export
	);

	altera_reset_sequencer #(
		.NUM_OUTPUTS                   (2),
		.ENABLE_DEASSERTION_INPUT_QUAL (0),
		.ENABLE_ASSERTION_SEQUENCE     (0),
		.ENABLE_DEASSERTION_SEQUENCE   (1),
		.MIN_ASRT_TIME                 (0),
		.ASRT_DELAY0                   (0),
		.DSRT_DELAY0                   (0),
		.ASRT_REMAP0                   (0),
		.DSRT_REMAP0                   (0),
		.DSRT_QUALCNT_0                (0),
		.ASRT_DELAY1                   (0),
		.DSRT_DELAY1                   (128),
		.ASRT_REMAP1                   (1),
		.DSRT_REMAP1                   (1),
		.DSRT_QUALCNT_1                (0),
		.ASRT_DELAY2                   (0),
		.DSRT_DELAY2                   (0),
		.ASRT_REMAP2                   (2),
		.DSRT_REMAP2                   (2),
		.DSRT_QUALCNT_2                (0),
		.ASRT_DELAY3                   (0),
		.DSRT_DELAY3                   (0),
		.ASRT_REMAP3                   (3),
		.DSRT_REMAP3                   (3),
		.DSRT_QUALCNT_3                (0),
		.ASRT_DELAY4                   (0),
		.DSRT_DELAY4                   (0),
		.ASRT_REMAP4                   (4),
		.DSRT_REMAP4                   (4),
		.DSRT_QUALCNT_4                (0),
		.ASRT_DELAY5                   (0),
		.DSRT_DELAY5                   (0),
		.ASRT_REMAP5                   (5),
		.DSRT_REMAP5                   (5),
		.DSRT_QUALCNT_5                (0),
		.ASRT_DELAY6                   (0),
		.DSRT_DELAY6                   (0),
		.ASRT_REMAP6                   (6),
		.DSRT_REMAP6                   (6),
		.DSRT_QUALCNT_6                (0),
		.ASRT_DELAY7                   (0),
		.DSRT_DELAY7                   (0),
		.ASRT_REMAP7                   (7),
		.DSRT_REMAP7                   (7),
		.DSRT_QUALCNT_7                (0),
		.ASRT_DELAY8                   (0),
		.DSRT_DELAY8                   (0),
		.ASRT_REMAP8                   (8),
		.DSRT_REMAP8                   (8),
		.DSRT_QUALCNT_8                (0),
		.ASRT_DELAY9                   (0),
		.DSRT_DELAY9                   (0),
		.ASRT_REMAP9                   (9),
		.DSRT_REMAP9                   (9),
		.DSRT_QUALCNT_9                (0),
		.ENABLE_CSR                    (0)
	) reset_sequencer_0 (
		.clk              (cpu_clk_out_clk),                    //        clk.clk
		.reset_in0        (~soc_reset_n),                       //  reset_in0.reset
		.reset_out0       (reset_sequencer_0_reset_out0_reset), // reset_out0.reset
		.reset_out1       (reset_sequencer_0_reset_out1_reset), // reset_out1.reset
		.reset_req_in0    (1'b0),                               // (terminated)
		.reset_in1        (1'b0),                               // (terminated)
		.reset_req_in1    (1'b0),                               // (terminated)
		.reset_in2        (1'b0),                               // (terminated)
		.reset_req_in2    (1'b0),                               // (terminated)
		.reset_in3        (1'b0),                               // (terminated)
		.reset_req_in3    (1'b0),                               // (terminated)
		.reset_in4        (1'b0),                               // (terminated)
		.reset_req_in4    (1'b0),                               // (terminated)
		.reset_in5        (1'b0),                               // (terminated)
		.reset_req_in5    (1'b0),                               // (terminated)
		.reset_in6        (1'b0),                               // (terminated)
		.reset_req_in6    (1'b0),                               // (terminated)
		.reset_in7        (1'b0),                               // (terminated)
		.reset_req_in7    (1'b0),                               // (terminated)
		.reset_in8        (1'b0),                               // (terminated)
		.reset_req_in8    (1'b0),                               // (terminated)
		.reset_in9        (1'b0),                               // (terminated)
		.reset_req_in9    (1'b0),                               // (terminated)
		.reset_req_out0   (),                                   // (terminated)
		.reset_req_out1   (),                                   // (terminated)
		.reset_out2       (),                                   // (terminated)
		.reset_req_out2   (),                                   // (terminated)
		.reset_out3       (),                                   // (terminated)
		.reset_req_out3   (),                                   // (terminated)
		.reset_out4       (),                                   // (terminated)
		.reset_req_out4   (),                                   // (terminated)
		.reset_out5       (),                                   // (terminated)
		.reset_req_out5   (),                                   // (terminated)
		.reset_out6       (),                                   // (terminated)
		.reset_req_out6   (),                                   // (terminated)
		.reset_out7       (),                                   // (terminated)
		.reset_req_out7   (),                                   // (terminated)
		.reset_out8       (),                                   // (terminated)
		.reset_req_out8   (),                                   // (terminated)
		.reset_out9       (),                                   // (terminated)
		.reset_req_out9   (),                                   // (terminated)
		.reset0_dsrt_qual (1'b0),                               // (terminated)
		.reset1_dsrt_qual (1'b0),                               // (terminated)
		.reset2_dsrt_qual (1'b0),                               // (terminated)
		.reset3_dsrt_qual (1'b0),                               // (terminated)
		.reset4_dsrt_qual (1'b0),                               // (terminated)
		.reset5_dsrt_qual (1'b0),                               // (terminated)
		.reset6_dsrt_qual (1'b0),                               // (terminated)
		.reset7_dsrt_qual (1'b0),                               // (terminated)
		.reset8_dsrt_qual (1'b0),                               // (terminated)
		.reset9_dsrt_qual (1'b0)                                // (terminated)
	);

	de10lite_sopc_sdram sdram (
		.clk            (pll_0_outclk1_clk),                        //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	de10lite_sopc_core_clk_freq soc_id (
		.clk      (cpu_clk_out_clk),                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_soc_id_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_soc_id_s1_readdata), //                    .readdata
		.in_port  (soc_id_export)                         // external_connection.export
	);

	de10lite_sopc_mm_interconnect_0 mm_interconnect_0 (
		.default_slave_axi_error_if_awid            (mm_interconnect_0_default_slave_axi_error_if_awid),    //           default_slave_axi_error_if.awid
		.default_slave_axi_error_if_awaddr          (mm_interconnect_0_default_slave_axi_error_if_awaddr),  //                                     .awaddr
		.default_slave_axi_error_if_awlen           (mm_interconnect_0_default_slave_axi_error_if_awlen),   //                                     .awlen
		.default_slave_axi_error_if_awsize          (mm_interconnect_0_default_slave_axi_error_if_awsize),  //                                     .awsize
		.default_slave_axi_error_if_awburst         (mm_interconnect_0_default_slave_axi_error_if_awburst), //                                     .awburst
		.default_slave_axi_error_if_awlock          (mm_interconnect_0_default_slave_axi_error_if_awlock),  //                                     .awlock
		.default_slave_axi_error_if_awcache         (mm_interconnect_0_default_slave_axi_error_if_awcache), //                                     .awcache
		.default_slave_axi_error_if_awprot          (mm_interconnect_0_default_slave_axi_error_if_awprot),  //                                     .awprot
		.default_slave_axi_error_if_awvalid         (mm_interconnect_0_default_slave_axi_error_if_awvalid), //                                     .awvalid
		.default_slave_axi_error_if_awready         (mm_interconnect_0_default_slave_axi_error_if_awready), //                                     .awready
		.default_slave_axi_error_if_wid             (mm_interconnect_0_default_slave_axi_error_if_wid),     //                                     .wid
		.default_slave_axi_error_if_wdata           (mm_interconnect_0_default_slave_axi_error_if_wdata),   //                                     .wdata
		.default_slave_axi_error_if_wstrb           (mm_interconnect_0_default_slave_axi_error_if_wstrb),   //                                     .wstrb
		.default_slave_axi_error_if_wlast           (mm_interconnect_0_default_slave_axi_error_if_wlast),   //                                     .wlast
		.default_slave_axi_error_if_wvalid          (mm_interconnect_0_default_slave_axi_error_if_wvalid),  //                                     .wvalid
		.default_slave_axi_error_if_wready          (mm_interconnect_0_default_slave_axi_error_if_wready),  //                                     .wready
		.default_slave_axi_error_if_bid             (mm_interconnect_0_default_slave_axi_error_if_bid),     //                                     .bid
		.default_slave_axi_error_if_bresp           (mm_interconnect_0_default_slave_axi_error_if_bresp),   //                                     .bresp
		.default_slave_axi_error_if_bvalid          (mm_interconnect_0_default_slave_axi_error_if_bvalid),  //                                     .bvalid
		.default_slave_axi_error_if_bready          (mm_interconnect_0_default_slave_axi_error_if_bready),  //                                     .bready
		.default_slave_axi_error_if_arid            (mm_interconnect_0_default_slave_axi_error_if_arid),    //                                     .arid
		.default_slave_axi_error_if_araddr          (mm_interconnect_0_default_slave_axi_error_if_araddr),  //                                     .araddr
		.default_slave_axi_error_if_arlen           (mm_interconnect_0_default_slave_axi_error_if_arlen),   //                                     .arlen
		.default_slave_axi_error_if_arsize          (mm_interconnect_0_default_slave_axi_error_if_arsize),  //                                     .arsize
		.default_slave_axi_error_if_arburst         (mm_interconnect_0_default_slave_axi_error_if_arburst), //                                     .arburst
		.default_slave_axi_error_if_arlock          (mm_interconnect_0_default_slave_axi_error_if_arlock),  //                                     .arlock
		.default_slave_axi_error_if_arcache         (mm_interconnect_0_default_slave_axi_error_if_arcache), //                                     .arcache
		.default_slave_axi_error_if_arprot          (mm_interconnect_0_default_slave_axi_error_if_arprot),  //                                     .arprot
		.default_slave_axi_error_if_arvalid         (mm_interconnect_0_default_slave_axi_error_if_arvalid), //                                     .arvalid
		.default_slave_axi_error_if_arready         (mm_interconnect_0_default_slave_axi_error_if_arready), //                                     .arready
		.default_slave_axi_error_if_rid             (mm_interconnect_0_default_slave_axi_error_if_rid),     //                                     .rid
		.default_slave_axi_error_if_rdata           (mm_interconnect_0_default_slave_axi_error_if_rdata),   //                                     .rdata
		.default_slave_axi_error_if_rresp           (mm_interconnect_0_default_slave_axi_error_if_rresp),   //                                     .rresp
		.default_slave_axi_error_if_rlast           (mm_interconnect_0_default_slave_axi_error_if_rlast),   //                                     .rlast
		.default_slave_axi_error_if_rvalid          (mm_interconnect_0_default_slave_axi_error_if_rvalid),  //                                     .rvalid
		.default_slave_axi_error_if_rready          (mm_interconnect_0_default_slave_axi_error_if_rready),  //                                     .rready
		.pll_0_outclk0_clk                          (cpu_clk_out_clk),                                      //                        pll_0_outclk0.clk
		.pll_0_outclk1_clk                          (pll_0_outclk1_clk),                                    //                        pll_0_outclk1.clk
		.avl_imem_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // avl_imem_reset_reset_bridge_in_reset.reset
		.sdram_reset_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                   //    sdram_reset_reset_bridge_in_reset.reset
		.avl_dmem_m0_address                        (avl_dmem_m0_address),                                  //                          avl_dmem_m0.address
		.avl_dmem_m0_waitrequest                    (avl_dmem_m0_waitrequest),                              //                                     .waitrequest
		.avl_dmem_m0_burstcount                     (avl_dmem_m0_burstcount),                               //                                     .burstcount
		.avl_dmem_m0_byteenable                     (avl_dmem_m0_byteenable),                               //                                     .byteenable
		.avl_dmem_m0_read                           (avl_dmem_m0_read),                                     //                                     .read
		.avl_dmem_m0_readdata                       (avl_dmem_m0_readdata),                                 //                                     .readdata
		.avl_dmem_m0_readdatavalid                  (avl_dmem_m0_readdatavalid),                            //                                     .readdatavalid
		.avl_dmem_m0_write                          (avl_dmem_m0_write),                                    //                                     .write
		.avl_dmem_m0_writedata                      (avl_dmem_m0_writedata),                                //                                     .writedata
		.avl_dmem_m0_debugaccess                    (avl_dmem_m0_debugaccess),                              //                                     .debugaccess
		.avl_dmem_m0_response                       (avl_dmem_m0_response),                                 //                                     .response
		.avl_imem_m0_address                        (avl_imem_m0_address),                                  //                          avl_imem_m0.address
		.avl_imem_m0_waitrequest                    (avl_imem_m0_waitrequest),                              //                                     .waitrequest
		.avl_imem_m0_burstcount                     (avl_imem_m0_burstcount),                               //                                     .burstcount
		.avl_imem_m0_byteenable                     (avl_imem_m0_byteenable),                               //                                     .byteenable
		.avl_imem_m0_read                           (avl_imem_m0_read),                                     //                                     .read
		.avl_imem_m0_readdata                       (avl_imem_m0_readdata),                                 //                                     .readdata
		.avl_imem_m0_readdatavalid                  (avl_imem_m0_readdatavalid),                            //                                     .readdatavalid
		.avl_imem_m0_write                          (avl_imem_m0_write),                                    //                                     .write
		.avl_imem_m0_writedata                      (avl_imem_m0_writedata),                                //                                     .writedata
		.avl_imem_m0_debugaccess                    (avl_imem_m0_debugaccess),                              //                                     .debugaccess
		.avl_imem_m0_response                       (avl_imem_m0_response),                                 //                                     .response
		.avl_uart_s0_address                        (mm_interconnect_0_avl_uart_s0_address),                //                          avl_uart_s0.address
		.avl_uart_s0_write                          (mm_interconnect_0_avl_uart_s0_write),                  //                                     .write
		.avl_uart_s0_read                           (mm_interconnect_0_avl_uart_s0_read),                   //                                     .read
		.avl_uart_s0_readdata                       (mm_interconnect_0_avl_uart_s0_readdata),               //                                     .readdata
		.avl_uart_s0_writedata                      (mm_interconnect_0_avl_uart_s0_writedata),              //                                     .writedata
		.avl_uart_s0_burstcount                     (mm_interconnect_0_avl_uart_s0_burstcount),             //                                     .burstcount
		.avl_uart_s0_byteenable                     (mm_interconnect_0_avl_uart_s0_byteenable),             //                                     .byteenable
		.avl_uart_s0_readdatavalid                  (mm_interconnect_0_avl_uart_s0_readdatavalid),          //                                     .readdatavalid
		.avl_uart_s0_waitrequest                    (mm_interconnect_0_avl_uart_s0_waitrequest),            //                                     .waitrequest
		.avl_uart_s0_debugaccess                    (mm_interconnect_0_avl_uart_s0_debugaccess),            //                                     .debugaccess
		.bld_id_s1_address                          (mm_interconnect_0_bld_id_s1_address),                  //                            bld_id_s1.address
		.bld_id_s1_readdata                         (mm_interconnect_0_bld_id_s1_readdata),                 //                                     .readdata
		.core_clk_freq_s1_address                   (mm_interconnect_0_core_clk_freq_s1_address),           //                     core_clk_freq_s1.address
		.core_clk_freq_s1_readdata                  (mm_interconnect_0_core_clk_freq_s1_readdata),          //                                     .readdata
		.onchip_ram_s1_address                      (mm_interconnect_0_onchip_ram_s1_address),              //                        onchip_ram_s1.address
		.onchip_ram_s1_write                        (mm_interconnect_0_onchip_ram_s1_write),                //                                     .write
		.onchip_ram_s1_readdata                     (mm_interconnect_0_onchip_ram_s1_readdata),             //                                     .readdata
		.onchip_ram_s1_writedata                    (mm_interconnect_0_onchip_ram_s1_writedata),            //                                     .writedata
		.onchip_ram_s1_byteenable                   (mm_interconnect_0_onchip_ram_s1_byteenable),           //                                     .byteenable
		.onchip_ram_s1_chipselect                   (mm_interconnect_0_onchip_ram_s1_chipselect),           //                                     .chipselect
		.onchip_ram_s1_clken                        (mm_interconnect_0_onchip_ram_s1_clken),                //                                     .clken
		.pio_led_s1_address                         (mm_interconnect_0_pio_led_s1_address),                 //                           pio_led_s1.address
		.pio_led_s1_write                           (mm_interconnect_0_pio_led_s1_write),                   //                                     .write
		.pio_led_s1_readdata                        (mm_interconnect_0_pio_led_s1_readdata),                //                                     .readdata
		.pio_led_s1_writedata                       (mm_interconnect_0_pio_led_s1_writedata),               //                                     .writedata
		.pio_led_s1_chipselect                      (mm_interconnect_0_pio_led_s1_chipselect),              //                                     .chipselect
		.pio_sw_s1_address                          (mm_interconnect_0_pio_sw_s1_address),                  //                            pio_sw_s1.address
		.pio_sw_s1_readdata                         (mm_interconnect_0_pio_sw_s1_readdata),                 //                                     .readdata
		.sdram_s1_address                           (mm_interconnect_0_sdram_s1_address),                   //                             sdram_s1.address
		.sdram_s1_write                             (mm_interconnect_0_sdram_s1_write),                     //                                     .write
		.sdram_s1_read                              (mm_interconnect_0_sdram_s1_read),                      //                                     .read
		.sdram_s1_readdata                          (mm_interconnect_0_sdram_s1_readdata),                  //                                     .readdata
		.sdram_s1_writedata                         (mm_interconnect_0_sdram_s1_writedata),                 //                                     .writedata
		.sdram_s1_byteenable                        (mm_interconnect_0_sdram_s1_byteenable),                //                                     .byteenable
		.sdram_s1_readdatavalid                     (mm_interconnect_0_sdram_s1_readdatavalid),             //                                     .readdatavalid
		.sdram_s1_waitrequest                       (mm_interconnect_0_sdram_s1_waitrequest),               //                                     .waitrequest
		.sdram_s1_chipselect                        (mm_interconnect_0_sdram_s1_chipselect),                //                                     .chipselect
		.soc_id_s1_address                          (mm_interconnect_0_soc_id_s1_address),                  //                            soc_id_s1.address
		.soc_id_s1_readdata                         (mm_interconnect_0_soc_id_s1_readdata)                  //                                     .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_sequencer_0_reset_out0_reset), // reset_in0.reset
		.clk            (cpu_clk_out_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (reset_sequencer_0_reset_out1_reset), // reset_in0.reset
		.clk            (cpu_clk_out_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (reset_sequencer_0_reset_out0_reset), // reset_in0.reset
		.clk            (pll_0_outclk1_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign cpu_rst_out_reset_n = ~rst_controller_001_reset_out_reset;

endmodule
